
module RAM(adress,datain,rw,enram,dataoutRAM); 

input enram;
input rw;
input [0:7] adress;
input [0:7] datain;
wire [0:255] selectList;
wire [0:2047] allResults;
output [0:7] dataoutRAM;

decoder d1(adress,enram,selectList); // 8x256 DECODER, SEND THE INPUTS

 genvar i;
  genvar j;
  
  generate

  for (i=0; i<256; i=i+1)  //LOOPS EVERY ADDRESS [0:255]
  begin : gen_loop
        for(j=0; j<8; j=j+1)  //LOOPS EVERY BIT [0:7]
        begin: gen_loop
        
			binaryCell bc1(datain[j],selectList[i],rw,allResults[(i*8)+j]);
			
        end
	
  end
  endgenerate
  
 //OR ALL BINARYCELL OUTPUTS 
assign dataoutRAM[0]=allResults[0]|allResults[8]|allResults[16]|allResults[24]|allResults[32]|allResults[40]|allResults[48]|allResults[56]|allResults[64]|allResults[72]|allResults[80]|allResults[88]|allResults[96]|allResults[104]|allResults[112]|allResults[120]|allResults[128]|allResults[136]|allResults[144]|allResults[152]|allResults[160]|allResults[168]|allResults[176]|allResults[184]|allResults[192]|allResults[200]|allResults[208]|allResults[216]|allResults[224]|allResults[232]|allResults[240]|allResults[248]|allResults[256]|allResults[264]|allResults[272]|allResults[280]|allResults[288]|allResults[296]|allResults[304]|allResults[312]|allResults[320]|allResults[328]|allResults[336]|allResults[344]|allResults[352]|allResults[360]|allResults[368]|allResults[376]|allResults[384]|allResults[392]|allResults[400]|allResults[408]|allResults[416]|allResults[424]|allResults[432]|allResults[440]|allResults[448]|allResults[456]|allResults[464]|allResults[472]|allResults[480]|allResults[488]|allResults[496]|allResults[504]|allResults[512]|allResults[520]|allResults[528]|allResults[536]|allResults[544]|allResults[552]|allResults[560]|allResults[568]|allResults[576]|allResults[584]|allResults[592]|allResults[600]|allResults[608]|allResults[616]|allResults[624]|allResults[632]|allResults[640]|allResults[648]|allResults[656]|allResults[664]|allResults[672]|allResults[680]|allResults[688]|allResults[696]|allResults[704]|allResults[712]|allResults[720]|allResults[728]|allResults[736]|allResults[744]|allResults[752]|allResults[760]|allResults[768]|allResults[776]|allResults[784]|allResults[792]|allResults[800]|allResults[808]|allResults[816]|allResults[824]|allResults[832]|allResults[840]|allResults[848]|allResults[856]|allResults[864]|allResults[872]|allResults[880]|allResults[888]|allResults[896]|allResults[904]|allResults[912]|allResults[920]|allResults[928]|allResults[936]|allResults[944]|allResults[952]|allResults[960]|allResults[968]|allResults[976]|allResults[984]|allResults[992]|allResults[1000]|allResults[1008]|allResults[1016]|allResults[1024]|allResults[1032]|allResults[1040]|allResults[1048]|allResults[1056]|allResults[1064]|allResults[1072]|allResults[1080]|allResults[1088]|allResults[1096]|allResults[1104]|allResults[1112]|allResults[1120]|allResults[1128]|allResults[1136]|allResults[1144]|allResults[1152]|allResults[1160]|allResults[1168]|allResults[1176]|allResults[1184]|allResults[1192]|allResults[1200]|allResults[1208]|allResults[1216]|allResults[1224]|allResults[1232]|allResults[1240]|allResults[1248]|allResults[1256]|allResults[1264]|allResults[1272]|allResults[1280]|allResults[1288]|allResults[1296]|allResults[1304]|allResults[1312]|allResults[1320]|allResults[1328]|allResults[1336]|allResults[1344]|allResults[1352]|allResults[1360]|allResults[1368]|allResults[1376]|allResults[1384]|allResults[1392]|allResults[1400]|allResults[1408]|allResults[1416]|allResults[1424]|allResults[1432]|allResults[1440]|allResults[1448]|allResults[1456]|allResults[1464]|allResults[1472]|allResults[1480]|allResults[1488]|allResults[1496]|allResults[1504]|allResults[1512]|allResults[1520]|allResults[1528]|allResults[1536]|allResults[1544]|allResults[1552]|allResults[1560]|allResults[1568]|allResults[1576]|allResults[1584]|allResults[1592]|allResults[1600]|allResults[1608]|allResults[1616]|allResults[1624]|allResults[1632]|allResults[1640]|allResults[1648]|allResults[1656]|allResults[1664]|allResults[1672]|allResults[1680]|allResults[1688]|allResults[1696]|allResults[1704]|allResults[1712]|allResults[1720]|allResults[1728]|allResults[1736]|allResults[1744]|allResults[1752]|allResults[1760]|allResults[1768]|allResults[1776]|allResults[1784]|allResults[1792]|allResults[1800]|allResults[1808]|allResults[1816]|allResults[1824]|allResults[1832]|allResults[1840]|allResults[1848]|allResults[1856]|allResults[1864]|allResults[1872]|allResults[1880]|allResults[1888]|allResults[1896]|allResults[1904]|allResults[1912]|allResults[1920]|allResults[1928]|allResults[1936]|allResults[1944]|allResults[1952]|allResults[1960]|allResults[1968]|allResults[1976]|allResults[1984]|allResults[1992]|allResults[2000]|allResults[2008]|allResults[2016]|allResults[2024]|allResults[2032]|allResults[2040];
assign dataoutRAM[1]=allResults[1]|allResults[9]|allResults[17]|allResults[25]|allResults[33]|allResults[41]|allResults[49]|allResults[57]|allResults[65]|allResults[73]|allResults[81]|allResults[89]|allResults[97]|allResults[105]|allResults[113]|allResults[121]|allResults[129]|allResults[137]|allResults[145]|allResults[153]|allResults[161]|allResults[169]|allResults[177]|allResults[185]|allResults[193]|allResults[201]|allResults[209]|allResults[217]|allResults[225]|allResults[233]|allResults[241]|allResults[249]|allResults[257]|allResults[265]|allResults[273]|allResults[281]|allResults[289]|allResults[297]|allResults[305]|allResults[313]|allResults[321]|allResults[329]|allResults[337]|allResults[345]|allResults[353]|allResults[361]|allResults[369]|allResults[377]|allResults[385]|allResults[393]|allResults[401]|allResults[409]|allResults[417]|allResults[425]|allResults[433]|allResults[441]|allResults[449]|allResults[457]|allResults[465]|allResults[473]|allResults[481]|allResults[489]|allResults[497]|allResults[505]|allResults[513]|allResults[521]|allResults[529]|allResults[537]|allResults[545]|allResults[553]|allResults[561]|allResults[569]|allResults[577]|allResults[585]|allResults[593]|allResults[601]|allResults[609]|allResults[617]|allResults[625]|allResults[633]|allResults[641]|allResults[649]|allResults[657]|allResults[665]|allResults[673]|allResults[681]|allResults[689]|allResults[697]|allResults[705]|allResults[713]|allResults[721]|allResults[729]|allResults[737]|allResults[745]|allResults[753]|allResults[761]|allResults[769]|allResults[777]|allResults[785]|allResults[793]|allResults[801]|allResults[809]|allResults[817]|allResults[825]|allResults[833]|allResults[841]|allResults[849]|allResults[857]|allResults[865]|allResults[873]|allResults[881]|allResults[889]|allResults[897]|allResults[905]|allResults[913]|allResults[921]|allResults[929]|allResults[937]|allResults[945]|allResults[953]|allResults[961]|allResults[969]|allResults[977]|allResults[985]|allResults[993]|allResults[1001]|allResults[1009]|allResults[1017]|allResults[1025]|allResults[1033]|allResults[1041]|allResults[1049]|allResults[1057]|allResults[1065]|allResults[1073]|allResults[1081]|allResults[1089]|allResults[1097]|allResults[1105]|allResults[1113]|allResults[1121]|allResults[1129]|allResults[1137]|allResults[1145]|allResults[1153]|allResults[1161]|allResults[1169]|allResults[1177]|allResults[1185]|allResults[1193]|allResults[1201]|allResults[1209]|allResults[1217]|allResults[1225]|allResults[1233]|allResults[1241]|allResults[1249]|allResults[1257]|allResults[1265]|allResults[1273]|allResults[1281]|allResults[1289]|allResults[1297]|allResults[1305]|allResults[1313]|allResults[1321]|allResults[1329]|allResults[1337]|allResults[1345]|allResults[1353]|allResults[1361]|allResults[1369]|allResults[1377]|allResults[1385]|allResults[1393]|allResults[1401]|allResults[1409]|allResults[1417]|allResults[1425]|allResults[1433]|allResults[1441]|allResults[1449]|allResults[1457]|allResults[1465]|allResults[1473]|allResults[1481]|allResults[1489]|allResults[1497]|allResults[1505]|allResults[1513]|allResults[1521]|allResults[1529]|allResults[1537]|allResults[1545]|allResults[1553]|allResults[1561]|allResults[1569]|allResults[1577]|allResults[1585]|allResults[1593]|allResults[1601]|allResults[1609]|allResults[1617]|allResults[1625]|allResults[1633]|allResults[1641]|allResults[1649]|allResults[1657]|allResults[1665]|allResults[1673]|allResults[1681]|allResults[1689]|allResults[1697]|allResults[1705]|allResults[1713]|allResults[1721]|allResults[1729]|allResults[1737]|allResults[1745]|allResults[1753]|allResults[1761]|allResults[1769]|allResults[1777]|allResults[1785]|allResults[1793]|allResults[1801]|allResults[1809]|allResults[1817]|allResults[1825]|allResults[1833]|allResults[1841]|allResults[1849]|allResults[1857]|allResults[1865]|allResults[1873]|allResults[1881]|allResults[1889]|allResults[1897]|allResults[1905]|allResults[1913]|allResults[1921]|allResults[1929]|allResults[1937]|allResults[1945]|allResults[1953]|allResults[1961]|allResults[1969]|allResults[1977]|allResults[1985]|allResults[1993]|allResults[2001]|allResults[2009]|allResults[2017]|allResults[2025]|allResults[2033]|allResults[2041];
assign dataoutRAM[2]=allResults[2]|allResults[10]|allResults[18]|allResults[26]|allResults[34]|allResults[42]|allResults[50]|allResults[58]|allResults[66]|allResults[74]|allResults[82]|allResults[90]|allResults[98]|allResults[106]|allResults[114]|allResults[122]|allResults[130]|allResults[138]|allResults[146]|allResults[154]|allResults[162]|allResults[170]|allResults[178]|allResults[186]|allResults[194]|allResults[202]|allResults[210]|allResults[218]|allResults[226]|allResults[234]|allResults[242]|allResults[250]|allResults[258]|allResults[266]|allResults[274]|allResults[282]|allResults[290]|allResults[298]|allResults[306]|allResults[314]|allResults[322]|allResults[330]|allResults[338]|allResults[346]|allResults[354]|allResults[362]|allResults[370]|allResults[378]|allResults[386]|allResults[394]|allResults[402]|allResults[410]|allResults[418]|allResults[426]|allResults[434]|allResults[442]|allResults[450]|allResults[458]|allResults[466]|allResults[474]|allResults[482]|allResults[490]|allResults[498]|allResults[506]|allResults[514]|allResults[522]|allResults[530]|allResults[538]|allResults[546]|allResults[554]|allResults[562]|allResults[570]|allResults[578]|allResults[586]|allResults[594]|allResults[602]|allResults[610]|allResults[618]|allResults[626]|allResults[634]|allResults[642]|allResults[650]|allResults[658]|allResults[666]|allResults[674]|allResults[682]|allResults[690]|allResults[698]|allResults[706]|allResults[714]|allResults[722]|allResults[730]|allResults[738]|allResults[746]|allResults[754]|allResults[762]|allResults[770]|allResults[778]|allResults[786]|allResults[794]|allResults[802]|allResults[810]|allResults[818]|allResults[826]|allResults[834]|allResults[842]|allResults[850]|allResults[858]|allResults[866]|allResults[874]|allResults[882]|allResults[890]|allResults[898]|allResults[906]|allResults[914]|allResults[922]|allResults[930]|allResults[938]|allResults[946]|allResults[954]|allResults[962]|allResults[970]|allResults[978]|allResults[986]|allResults[994]|allResults[1002]|allResults[1010]|allResults[1018]|allResults[1026]|allResults[1034]|allResults[1042]|allResults[1050]|allResults[1058]|allResults[1066]|allResults[1074]|allResults[1082]|allResults[1090]|allResults[1098]|allResults[1106]|allResults[1114]|allResults[1122]|allResults[1130]|allResults[1138]|allResults[1146]|allResults[1154]|allResults[1162]|allResults[1170]|allResults[1178]|allResults[1186]|allResults[1194]|allResults[1202]|allResults[1210]|allResults[1218]|allResults[1226]|allResults[1234]|allResults[1242]|allResults[1250]|allResults[1258]|allResults[1266]|allResults[1274]|allResults[1282]|allResults[1290]|allResults[1298]|allResults[1306]|allResults[1314]|allResults[1322]|allResults[1330]|allResults[1338]|allResults[1346]|allResults[1354]|allResults[1362]|allResults[1370]|allResults[1378]|allResults[1386]|allResults[1394]|allResults[1402]|allResults[1410]|allResults[1418]|allResults[1426]|allResults[1434]|allResults[1442]|allResults[1450]|allResults[1458]|allResults[1466]|allResults[1474]|allResults[1482]|allResults[1490]|allResults[1498]|allResults[1506]|allResults[1514]|allResults[1522]|allResults[1530]|allResults[1538]|allResults[1546]|allResults[1554]|allResults[1562]|allResults[1570]|allResults[1578]|allResults[1586]|allResults[1594]|allResults[1602]|allResults[1610]|allResults[1618]|allResults[1626]|allResults[1634]|allResults[1642]|allResults[1650]|allResults[1658]|allResults[1666]|allResults[1674]|allResults[1682]|allResults[1690]|allResults[1698]|allResults[1706]|allResults[1714]|allResults[1722]|allResults[1730]|allResults[1738]|allResults[1746]|allResults[1754]|allResults[1762]|allResults[1770]|allResults[1778]|allResults[1786]|allResults[1794]|allResults[1802]|allResults[1810]|allResults[1818]|allResults[1826]|allResults[1834]|allResults[1842]|allResults[1850]|allResults[1858]|allResults[1866]|allResults[1874]|allResults[1882]|allResults[1890]|allResults[1898]|allResults[1906]|allResults[1914]|allResults[1922]|allResults[1930]|allResults[1938]|allResults[1946]|allResults[1954]|allResults[1962]|allResults[1970]|allResults[1978]|allResults[1986]|allResults[1994]|allResults[2002]|allResults[2010]|allResults[2018]|allResults[2026]|allResults[2034]|allResults[2042];
assign dataoutRAM[3]=allResults[3]|allResults[11]|allResults[19]|allResults[27]|allResults[35]|allResults[43]|allResults[51]|allResults[59]|allResults[67]|allResults[75]|allResults[83]|allResults[91]|allResults[99]|allResults[107]|allResults[115]|allResults[123]|allResults[131]|allResults[139]|allResults[147]|allResults[155]|allResults[163]|allResults[171]|allResults[179]|allResults[187]|allResults[195]|allResults[203]|allResults[211]|allResults[219]|allResults[227]|allResults[235]|allResults[243]|allResults[251]|allResults[259]|allResults[267]|allResults[275]|allResults[283]|allResults[291]|allResults[299]|allResults[307]|allResults[315]|allResults[323]|allResults[331]|allResults[339]|allResults[347]|allResults[355]|allResults[363]|allResults[371]|allResults[379]|allResults[387]|allResults[395]|allResults[403]|allResults[411]|allResults[419]|allResults[427]|allResults[435]|allResults[443]|allResults[451]|allResults[459]|allResults[467]|allResults[475]|allResults[483]|allResults[491]|allResults[499]|allResults[507]|allResults[515]|allResults[523]|allResults[531]|allResults[539]|allResults[547]|allResults[555]|allResults[563]|allResults[571]|allResults[579]|allResults[587]|allResults[595]|allResults[603]|allResults[611]|allResults[619]|allResults[627]|allResults[635]|allResults[643]|allResults[651]|allResults[659]|allResults[667]|allResults[675]|allResults[683]|allResults[691]|allResults[699]|allResults[707]|allResults[715]|allResults[723]|allResults[731]|allResults[739]|allResults[747]|allResults[755]|allResults[763]|allResults[771]|allResults[779]|allResults[787]|allResults[795]|allResults[803]|allResults[811]|allResults[819]|allResults[827]|allResults[835]|allResults[843]|allResults[851]|allResults[859]|allResults[867]|allResults[875]|allResults[883]|allResults[891]|allResults[899]|allResults[907]|allResults[915]|allResults[923]|allResults[931]|allResults[939]|allResults[947]|allResults[955]|allResults[963]|allResults[971]|allResults[979]|allResults[987]|allResults[995]|allResults[1003]|allResults[1011]|allResults[1019]|allResults[1027]|allResults[1035]|allResults[1043]|allResults[1051]|allResults[1059]|allResults[1067]|allResults[1075]|allResults[1083]|allResults[1091]|allResults[1099]|allResults[1107]|allResults[1115]|allResults[1123]|allResults[1131]|allResults[1139]|allResults[1147]|allResults[1155]|allResults[1163]|allResults[1171]|allResults[1179]|allResults[1187]|allResults[1195]|allResults[1203]|allResults[1211]|allResults[1219]|allResults[1227]|allResults[1235]|allResults[1243]|allResults[1251]|allResults[1259]|allResults[1267]|allResults[1275]|allResults[1283]|allResults[1291]|allResults[1299]|allResults[1307]|allResults[1315]|allResults[1323]|allResults[1331]|allResults[1339]|allResults[1347]|allResults[1355]|allResults[1363]|allResults[1371]|allResults[1379]|allResults[1387]|allResults[1395]|allResults[1403]|allResults[1411]|allResults[1419]|allResults[1427]|allResults[1435]|allResults[1443]|allResults[1451]|allResults[1459]|allResults[1467]|allResults[1475]|allResults[1483]|allResults[1491]|allResults[1499]|allResults[1507]|allResults[1515]|allResults[1523]|allResults[1531]|allResults[1539]|allResults[1547]|allResults[1555]|allResults[1563]|allResults[1571]|allResults[1579]|allResults[1587]|allResults[1595]|allResults[1603]|allResults[1611]|allResults[1619]|allResults[1627]|allResults[1635]|allResults[1643]|allResults[1651]|allResults[1659]|allResults[1667]|allResults[1675]|allResults[1683]|allResults[1691]|allResults[1699]|allResults[1707]|allResults[1715]|allResults[1723]|allResults[1731]|allResults[1739]|allResults[1747]|allResults[1755]|allResults[1763]|allResults[1771]|allResults[1779]|allResults[1787]|allResults[1795]|allResults[1803]|allResults[1811]|allResults[1819]|allResults[1827]|allResults[1835]|allResults[1843]|allResults[1851]|allResults[1859]|allResults[1867]|allResults[1875]|allResults[1883]|allResults[1891]|allResults[1899]|allResults[1907]|allResults[1915]|allResults[1923]|allResults[1931]|allResults[1939]|allResults[1947]|allResults[1955]|allResults[1963]|allResults[1971]|allResults[1979]|allResults[1987]|allResults[1995]|allResults[2003]|allResults[2011]|allResults[2019]|allResults[2027]|allResults[2035]|allResults[2043];
assign dataoutRAM[4]=allResults[4]|allResults[12]|allResults[20]|allResults[28]|allResults[36]|allResults[44]|allResults[52]|allResults[60]|allResults[68]|allResults[76]|allResults[84]|allResults[92]|allResults[100]|allResults[108]|allResults[116]|allResults[124]|allResults[132]|allResults[140]|allResults[148]|allResults[156]|allResults[164]|allResults[172]|allResults[180]|allResults[188]|allResults[196]|allResults[204]|allResults[212]|allResults[220]|allResults[228]|allResults[236]|allResults[244]|allResults[252]|allResults[260]|allResults[268]|allResults[276]|allResults[284]|allResults[292]|allResults[300]|allResults[308]|allResults[316]|allResults[324]|allResults[332]|allResults[340]|allResults[348]|allResults[356]|allResults[364]|allResults[372]|allResults[380]|allResults[388]|allResults[396]|allResults[404]|allResults[412]|allResults[420]|allResults[428]|allResults[436]|allResults[444]|allResults[452]|allResults[460]|allResults[468]|allResults[476]|allResults[484]|allResults[492]|allResults[500]|allResults[508]|allResults[516]|allResults[524]|allResults[532]|allResults[540]|allResults[548]|allResults[556]|allResults[564]|allResults[572]|allResults[580]|allResults[588]|allResults[596]|allResults[604]|allResults[612]|allResults[620]|allResults[628]|allResults[636]|allResults[644]|allResults[652]|allResults[660]|allResults[668]|allResults[676]|allResults[684]|allResults[692]|allResults[700]|allResults[708]|allResults[716]|allResults[724]|allResults[732]|allResults[740]|allResults[748]|allResults[756]|allResults[764]|allResults[772]|allResults[780]|allResults[788]|allResults[796]|allResults[804]|allResults[812]|allResults[820]|allResults[828]|allResults[836]|allResults[844]|allResults[852]|allResults[860]|allResults[868]|allResults[876]|allResults[884]|allResults[892]|allResults[900]|allResults[908]|allResults[916]|allResults[924]|allResults[932]|allResults[940]|allResults[948]|allResults[956]|allResults[964]|allResults[972]|allResults[980]|allResults[988]|allResults[996]|allResults[1004]|allResults[1012]|allResults[1020]|allResults[1028]|allResults[1036]|allResults[1044]|allResults[1052]|allResults[1060]|allResults[1068]|allResults[1076]|allResults[1084]|allResults[1092]|allResults[1100]|allResults[1108]|allResults[1116]|allResults[1124]|allResults[1132]|allResults[1140]|allResults[1148]|allResults[1156]|allResults[1164]|allResults[1172]|allResults[1180]|allResults[1188]|allResults[1196]|allResults[1204]|allResults[1212]|allResults[1220]|allResults[1228]|allResults[1236]|allResults[1244]|allResults[1252]|allResults[1260]|allResults[1268]|allResults[1276]|allResults[1284]|allResults[1292]|allResults[1300]|allResults[1308]|allResults[1316]|allResults[1324]|allResults[1332]|allResults[1340]|allResults[1348]|allResults[1356]|allResults[1364]|allResults[1372]|allResults[1380]|allResults[1388]|allResults[1396]|allResults[1404]|allResults[1412]|allResults[1420]|allResults[1428]|allResults[1436]|allResults[1444]|allResults[1452]|allResults[1460]|allResults[1468]|allResults[1476]|allResults[1484]|allResults[1492]|allResults[1500]|allResults[1508]|allResults[1516]|allResults[1524]|allResults[1532]|allResults[1540]|allResults[1548]|allResults[1556]|allResults[1564]|allResults[1572]|allResults[1580]|allResults[1588]|allResults[1596]|allResults[1604]|allResults[1612]|allResults[1620]|allResults[1628]|allResults[1636]|allResults[1644]|allResults[1652]|allResults[1660]|allResults[1668]|allResults[1676]|allResults[1684]|allResults[1692]|allResults[1700]|allResults[1708]|allResults[1716]|allResults[1724]|allResults[1732]|allResults[1740]|allResults[1748]|allResults[1756]|allResults[1764]|allResults[1772]|allResults[1780]|allResults[1788]|allResults[1796]|allResults[1804]|allResults[1812]|allResults[1820]|allResults[1828]|allResults[1836]|allResults[1844]|allResults[1852]|allResults[1860]|allResults[1868]|allResults[1876]|allResults[1884]|allResults[1892]|allResults[1900]|allResults[1908]|allResults[1916]|allResults[1924]|allResults[1932]|allResults[1940]|allResults[1948]|allResults[1956]|allResults[1964]|allResults[1972]|allResults[1980]|allResults[1988]|allResults[1996]|allResults[2004]|allResults[2012]|allResults[2020]|allResults[2028]|allResults[2036]|allResults[2044];
assign dataoutRAM[5]=allResults[5]|allResults[13]|allResults[21]|allResults[29]|allResults[37]|allResults[45]|allResults[53]|allResults[61]|allResults[69]|allResults[77]|allResults[85]|allResults[93]|allResults[101]|allResults[109]|allResults[117]|allResults[125]|allResults[133]|allResults[141]|allResults[149]|allResults[157]|allResults[165]|allResults[173]|allResults[181]|allResults[189]|allResults[197]|allResults[205]|allResults[213]|allResults[221]|allResults[229]|allResults[237]|allResults[245]|allResults[253]|allResults[261]|allResults[269]|allResults[277]|allResults[285]|allResults[293]|allResults[301]|allResults[309]|allResults[317]|allResults[325]|allResults[333]|allResults[341]|allResults[349]|allResults[357]|allResults[365]|allResults[373]|allResults[381]|allResults[389]|allResults[397]|allResults[405]|allResults[413]|allResults[421]|allResults[429]|allResults[437]|allResults[445]|allResults[453]|allResults[461]|allResults[469]|allResults[477]|allResults[485]|allResults[493]|allResults[501]|allResults[509]|allResults[517]|allResults[525]|allResults[533]|allResults[541]|allResults[549]|allResults[557]|allResults[565]|allResults[573]|allResults[581]|allResults[589]|allResults[597]|allResults[605]|allResults[613]|allResults[621]|allResults[629]|allResults[637]|allResults[645]|allResults[653]|allResults[661]|allResults[669]|allResults[677]|allResults[685]|allResults[693]|allResults[701]|allResults[709]|allResults[717]|allResults[725]|allResults[733]|allResults[741]|allResults[749]|allResults[757]|allResults[765]|allResults[773]|allResults[781]|allResults[789]|allResults[797]|allResults[805]|allResults[813]|allResults[821]|allResults[829]|allResults[837]|allResults[845]|allResults[853]|allResults[861]|allResults[869]|allResults[877]|allResults[885]|allResults[893]|allResults[901]|allResults[909]|allResults[917]|allResults[925]|allResults[933]|allResults[941]|allResults[949]|allResults[957]|allResults[965]|allResults[973]|allResults[981]|allResults[989]|allResults[997]|allResults[1005]|allResults[1013]|allResults[1021]|allResults[1029]|allResults[1037]|allResults[1045]|allResults[1053]|allResults[1061]|allResults[1069]|allResults[1077]|allResults[1085]|allResults[1093]|allResults[1101]|allResults[1109]|allResults[1117]|allResults[1125]|allResults[1133]|allResults[1141]|allResults[1149]|allResults[1157]|allResults[1165]|allResults[1173]|allResults[1181]|allResults[1189]|allResults[1197]|allResults[1205]|allResults[1213]|allResults[1221]|allResults[1229]|allResults[1237]|allResults[1245]|allResults[1253]|allResults[1261]|allResults[1269]|allResults[1277]|allResults[1285]|allResults[1293]|allResults[1301]|allResults[1309]|allResults[1317]|allResults[1325]|allResults[1333]|allResults[1341]|allResults[1349]|allResults[1357]|allResults[1365]|allResults[1373]|allResults[1381]|allResults[1389]|allResults[1397]|allResults[1405]|allResults[1413]|allResults[1421]|allResults[1429]|allResults[1437]|allResults[1445]|allResults[1453]|allResults[1461]|allResults[1469]|allResults[1477]|allResults[1485]|allResults[1493]|allResults[1501]|allResults[1509]|allResults[1517]|allResults[1525]|allResults[1533]|allResults[1541]|allResults[1549]|allResults[1557]|allResults[1565]|allResults[1573]|allResults[1581]|allResults[1589]|allResults[1597]|allResults[1605]|allResults[1613]|allResults[1621]|allResults[1629]|allResults[1637]|allResults[1645]|allResults[1653]|allResults[1661]|allResults[1669]|allResults[1677]|allResults[1685]|allResults[1693]|allResults[1701]|allResults[1709]|allResults[1717]|allResults[1725]|allResults[1733]|allResults[1741]|allResults[1749]|allResults[1757]|allResults[1765]|allResults[1773]|allResults[1781]|allResults[1789]|allResults[1797]|allResults[1805]|allResults[1813]|allResults[1821]|allResults[1829]|allResults[1837]|allResults[1845]|allResults[1853]|allResults[1861]|allResults[1869]|allResults[1877]|allResults[1885]|allResults[1893]|allResults[1901]|allResults[1909]|allResults[1917]|allResults[1925]|allResults[1933]|allResults[1941]|allResults[1949]|allResults[1957]|allResults[1965]|allResults[1973]|allResults[1981]|allResults[1989]|allResults[1997]|allResults[2005]|allResults[2013]|allResults[2021]|allResults[2029]|allResults[2037]|allResults[2045];
assign dataoutRAM[6]=allResults[6]|allResults[14]|allResults[22]|allResults[30]|allResults[38]|allResults[46]|allResults[54]|allResults[62]|allResults[70]|allResults[78]|allResults[86]|allResults[94]|allResults[102]|allResults[110]|allResults[118]|allResults[126]|allResults[134]|allResults[142]|allResults[150]|allResults[158]|allResults[166]|allResults[174]|allResults[182]|allResults[190]|allResults[198]|allResults[206]|allResults[214]|allResults[222]|allResults[230]|allResults[238]|allResults[246]|allResults[254]|allResults[262]|allResults[270]|allResults[278]|allResults[286]|allResults[294]|allResults[302]|allResults[310]|allResults[318]|allResults[326]|allResults[334]|allResults[342]|allResults[350]|allResults[358]|allResults[366]|allResults[374]|allResults[382]|allResults[390]|allResults[398]|allResults[406]|allResults[414]|allResults[422]|allResults[430]|allResults[438]|allResults[446]|allResults[454]|allResults[462]|allResults[470]|allResults[478]|allResults[486]|allResults[494]|allResults[502]|allResults[510]|allResults[518]|allResults[526]|allResults[534]|allResults[542]|allResults[550]|allResults[558]|allResults[566]|allResults[574]|allResults[582]|allResults[590]|allResults[598]|allResults[606]|allResults[614]|allResults[622]|allResults[630]|allResults[638]|allResults[646]|allResults[654]|allResults[662]|allResults[670]|allResults[678]|allResults[686]|allResults[694]|allResults[702]|allResults[710]|allResults[718]|allResults[726]|allResults[734]|allResults[742]|allResults[750]|allResults[758]|allResults[766]|allResults[774]|allResults[782]|allResults[790]|allResults[798]|allResults[806]|allResults[814]|allResults[822]|allResults[830]|allResults[838]|allResults[846]|allResults[854]|allResults[862]|allResults[870]|allResults[878]|allResults[886]|allResults[894]|allResults[902]|allResults[910]|allResults[918]|allResults[926]|allResults[934]|allResults[942]|allResults[950]|allResults[958]|allResults[966]|allResults[974]|allResults[982]|allResults[990]|allResults[998]|allResults[1006]|allResults[1014]|allResults[1022]|allResults[1030]|allResults[1038]|allResults[1046]|allResults[1054]|allResults[1062]|allResults[1070]|allResults[1078]|allResults[1086]|allResults[1094]|allResults[1102]|allResults[1110]|allResults[1118]|allResults[1126]|allResults[1134]|allResults[1142]|allResults[1150]|allResults[1158]|allResults[1166]|allResults[1174]|allResults[1182]|allResults[1190]|allResults[1198]|allResults[1206]|allResults[1214]|allResults[1222]|allResults[1230]|allResults[1238]|allResults[1246]|allResults[1254]|allResults[1262]|allResults[1270]|allResults[1278]|allResults[1286]|allResults[1294]|allResults[1302]|allResults[1310]|allResults[1318]|allResults[1326]|allResults[1334]|allResults[1342]|allResults[1350]|allResults[1358]|allResults[1366]|allResults[1374]|allResults[1382]|allResults[1390]|allResults[1398]|allResults[1406]|allResults[1414]|allResults[1422]|allResults[1430]|allResults[1438]|allResults[1446]|allResults[1454]|allResults[1462]|allResults[1470]|allResults[1478]|allResults[1486]|allResults[1494]|allResults[1502]|allResults[1510]|allResults[1518]|allResults[1526]|allResults[1534]|allResults[1542]|allResults[1550]|allResults[1558]|allResults[1566]|allResults[1574]|allResults[1582]|allResults[1590]|allResults[1598]|allResults[1606]|allResults[1614]|allResults[1622]|allResults[1630]|allResults[1638]|allResults[1646]|allResults[1654]|allResults[1662]|allResults[1670]|allResults[1678]|allResults[1686]|allResults[1694]|allResults[1702]|allResults[1710]|allResults[1718]|allResults[1726]|allResults[1734]|allResults[1742]|allResults[1750]|allResults[1758]|allResults[1766]|allResults[1774]|allResults[1782]|allResults[1790]|allResults[1798]|allResults[1806]|allResults[1814]|allResults[1822]|allResults[1830]|allResults[1838]|allResults[1846]|allResults[1854]|allResults[1862]|allResults[1870]|allResults[1878]|allResults[1886]|allResults[1894]|allResults[1902]|allResults[1910]|allResults[1918]|allResults[1926]|allResults[1934]|allResults[1942]|allResults[1950]|allResults[1958]|allResults[1966]|allResults[1974]|allResults[1982]|allResults[1990]|allResults[1998]|allResults[2006]|allResults[2014]|allResults[2022]|allResults[2030]|allResults[2038]|allResults[2046];
assign dataoutRAM[7]=allResults[7]|allResults[15]|allResults[23]|allResults[31]|allResults[39]|allResults[47]|allResults[55]|allResults[63]|allResults[71]|allResults[79]|allResults[87]|allResults[95]|allResults[103]|allResults[111]|allResults[119]|allResults[127]|allResults[135]|allResults[143]|allResults[151]|allResults[159]|allResults[167]|allResults[175]|allResults[183]|allResults[191]|allResults[199]|allResults[207]|allResults[215]|allResults[223]|allResults[231]|allResults[239]|allResults[247]|allResults[255]|allResults[263]|allResults[271]|allResults[279]|allResults[287]|allResults[295]|allResults[303]|allResults[311]|allResults[319]|allResults[327]|allResults[335]|allResults[343]|allResults[351]|allResults[359]|allResults[367]|allResults[375]|allResults[383]|allResults[391]|allResults[399]|allResults[407]|allResults[415]|allResults[423]|allResults[431]|allResults[439]|allResults[447]|allResults[455]|allResults[463]|allResults[471]|allResults[479]|allResults[487]|allResults[495]|allResults[503]|allResults[511]|allResults[519]|allResults[527]|allResults[535]|allResults[543]|allResults[551]|allResults[559]|allResults[567]|allResults[575]|allResults[583]|allResults[591]|allResults[599]|allResults[607]|allResults[615]|allResults[623]|allResults[631]|allResults[639]|allResults[647]|allResults[655]|allResults[663]|allResults[671]|allResults[679]|allResults[687]|allResults[695]|allResults[703]|allResults[711]|allResults[719]|allResults[727]|allResults[735]|allResults[743]|allResults[751]|allResults[759]|allResults[767]|allResults[775]|allResults[783]|allResults[791]|allResults[799]|allResults[807]|allResults[815]|allResults[823]|allResults[831]|allResults[839]|allResults[847]|allResults[855]|allResults[863]|allResults[871]|allResults[879]|allResults[887]|allResults[895]|allResults[903]|allResults[911]|allResults[919]|allResults[927]|allResults[935]|allResults[943]|allResults[951]|allResults[959]|allResults[967]|allResults[975]|allResults[983]|allResults[991]|allResults[999]|allResults[1007]|allResults[1015]|allResults[1023]|allResults[1031]|allResults[1039]|allResults[1047]|allResults[1055]|allResults[1063]|allResults[1071]|allResults[1079]|allResults[1087]|allResults[1095]|allResults[1103]|allResults[1111]|allResults[1119]|allResults[1127]|allResults[1135]|allResults[1143]|allResults[1151]|allResults[1159]|allResults[1167]|allResults[1175]|allResults[1183]|allResults[1191]|allResults[1199]|allResults[1207]|allResults[1215]|allResults[1223]|allResults[1231]|allResults[1239]|allResults[1247]|allResults[1255]|allResults[1263]|allResults[1271]|allResults[1279]|allResults[1287]|allResults[1295]|allResults[1303]|allResults[1311]|allResults[1319]|allResults[1327]|allResults[1335]|allResults[1343]|allResults[1351]|allResults[1359]|allResults[1367]|allResults[1375]|allResults[1383]|allResults[1391]|allResults[1399]|allResults[1407]|allResults[1415]|allResults[1423]|allResults[1431]|allResults[1439]|allResults[1447]|allResults[1455]|allResults[1463]|allResults[1471]|allResults[1479]|allResults[1487]|allResults[1495]|allResults[1503]|allResults[1511]|allResults[1519]|allResults[1527]|allResults[1535]|allResults[1543]|allResults[1551]|allResults[1559]|allResults[1567]|allResults[1575]|allResults[1583]|allResults[1591]|allResults[1599]|allResults[1607]|allResults[1615]|allResults[1623]|allResults[1631]|allResults[1639]|allResults[1647]|allResults[1655]|allResults[1663]|allResults[1671]|allResults[1679]|allResults[1687]|allResults[1695]|allResults[1703]|allResults[1711]|allResults[1719]|allResults[1727]|allResults[1735]|allResults[1743]|allResults[1751]|allResults[1759]|allResults[1767]|allResults[1775]|allResults[1783]|allResults[1791]|allResults[1799]|allResults[1807]|allResults[1815]|allResults[1823]|allResults[1831]|allResults[1839]|allResults[1847]|allResults[1855]|allResults[1863]|allResults[1871]|allResults[1879]|allResults[1887]|allResults[1895]|allResults[1903]|allResults[1911]|allResults[1919]|allResults[1927]|allResults[1935]|allResults[1943]|allResults[1951]|allResults[1959]|allResults[1967]|allResults[1975]|allResults[1983]|allResults[1991]|allResults[1999]|allResults[2007]|allResults[2015]|allResults[2023]|allResults[2031]|allResults[2039]|allResults[2047];


endmodule




