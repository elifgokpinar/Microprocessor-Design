module ROM(addr,enrom,data);
input [0:7] addr;
input enrom;
output reg [0:12] data; 
always@ (*)
begin
	 if(enrom)
	 begin
	   case(addr)
			8'b00000000 : data = 13'b0000011110000;
			8'b00000001 : data = 13'b0000011110000; //Literal type ADD
			8'b00000010 : data = 13'b0111100000000; //Register type STORE
			8'b00000011 : data = 13'b0100000000000; //Register type ADD
			8'b00000100 : data = 13'b0100000000000; 
			8'b00000101 : data = 13'b0000000000101;
			8'b00000110 : data = 13'b0000000000110;
			8'b00000111 : data = 13'b0000000000111;
			8'b00001000 : data = 13'b0000000001000;
			8'b00001001 : data = 13'b0000000001001;
			8'b00001010 : data = 13'b0000000001010;
			8'b00001011 : data = 13'b0000000001011;
			8'b00001100 : data = 13'b0000000001100;
			8'b00001101 : data = 13'b0000000001101;
			8'b00001110 : data = 13'b0000000001110;
			8'b00001111 : data = 13'b0000000001111;
			8'b00010000 : data = 13'b0000000010000;
			8'b00010001 : data = 13'b0000000010001;
			8'b00010010 : data = 13'b0000000010010;
			8'b00010011 : data = 13'b0000000010011;
			8'b00010100 : data = 13'b0000000010100;
			8'b00010101 : data = 13'b0000000010101;
			8'b00010110 : data = 13'b0000000010110;
			8'b00010111 : data = 13'b0000000010111;
			8'b00011000 : data = 13'b0000000011000;
			8'b00011001 : data = 13'b0000000011001;
			8'b00011010 : data = 13'b0000000011010;
			8'b00011011 : data = 13'b0000000011011;
			8'b00011100 : data = 13'b0000000011100;
			8'b00011101 : data = 13'b0000000011101;
			8'b00011110 : data = 13'b0000000011110;
			8'b00011111 : data = 13'b0000000011111;
			8'b00100000 : data = 13'b0000000100000;
			8'b00100001 : data = 13'b0000000100001;
			8'b00100010 : data = 13'b0000000100010;
			8'b00100011 : data = 13'b0000000100011;
			8'b00100100 : data = 13'b0000000100100;
			8'b00100101 : data = 13'b0000000100101;
			8'b00100110 : data = 13'b0000000100110;
			8'b00100111 : data = 13'b0000000100111;
			8'b00101000 : data = 13'b0000000101000;
			8'b00101001 : data = 13'b0000000101001;
			8'b00101010 : data = 13'b0000000101010;
			8'b00101011 : data = 13'b0000000101011;
			8'b00101100 : data = 13'b0000000101100;
			8'b00101101 : data = 13'b0000000101101;
			8'b00101110 : data = 13'b0000000101110;
			8'b00101111 : data = 13'b0000000101111;
			8'b00110000 : data = 13'b0000000110000;
			8'b00110001 : data = 13'b0000000110001;
			8'b00110010 : data = 13'b0000000110010;
			8'b00110011 : data = 13'b0000000110011;
			8'b00110100 : data = 13'b0000000110100;
			8'b00110101 : data = 13'b0000000110101;
			8'b00110110 : data = 13'b0000000110110;
			8'b00110111 : data = 13'b0000000110111;
			8'b00111000 : data = 13'b0000000111000;
			8'b00111001 : data = 13'b0000000111001;
			8'b00111010 : data = 13'b0000000111010;
			8'b00111011 : data = 13'b0000000111011;
			8'b00111100 : data = 13'b0000000111100;
			8'b00111101 : data = 13'b0000000111101;
			8'b00111110 : data = 13'b0000000111110;
			8'b00111111 : data = 13'b0000000111111;
			8'b01000000 : data = 13'b0000001000000;
			8'b01000001 : data = 13'b0000001000001;
			8'b01000010 : data = 13'b0000001000010;
			8'b01000011 : data = 13'b0000001000011;
			8'b01000100 : data = 13'b0000001000100;
			8'b01000101 : data = 13'b0000001000101;
			8'b01000110 : data = 13'b0000001000110;
			8'b01000111 : data = 13'b0000001000111;
			8'b01001000 : data = 13'b0000001001000;
			8'b01001001 : data = 13'b0000001001001;
			8'b01001010 : data = 13'b0000001001010;
			8'b01001011 : data = 13'b0000001001011;
			8'b01001100 : data = 13'b0000001001100;
			8'b01001101 : data = 13'b0000001001101;
			8'b01001110 : data = 13'b0000001001110;
			8'b01001111 : data = 13'b0000001001111;
			8'b01010000 : data = 13'b0000001010000;
			8'b01010001 : data = 13'b0000001010001;
			8'b01010010 : data = 13'b0000001010010;
			8'b01010011 : data = 13'b0000001010011;
			8'b01010100 : data = 13'b0000001010100;
			8'b01010101 : data = 13'b0000001010101;
			8'b01010110 : data = 13'b0000001010110;
			8'b01010111 : data = 13'b0000001010111;
			8'b01011000 : data = 13'b0000001011000;
			8'b01011001 : data = 13'b0000001011001;
			8'b01011010 : data = 13'b0000001011010;
			8'b01011011 : data = 13'b0000001011011;
			8'b01011100 : data = 13'b0000001011100;
			8'b01011101 : data = 13'b0000001011101;
			8'b01011110 : data = 13'b0000001011110;
			8'b01011111 : data = 13'b0000001011111;
			8'b01100000 : data = 13'b0000001100000;
			8'b01100001 : data = 13'b0000001100001;
			8'b01100010 : data = 13'b0000001100010;
			8'b01100011 : data = 13'b0000001100011;
			8'b01100100 : data = 13'b0000001100100;
			8'b01100101 : data = 13'b0000001100101;
			8'b01100110 : data = 13'b0000001100110;
			8'b01100111 : data = 13'b0000001100111;
			8'b01101000 : data = 13'b0000001101000;
			8'b01101001 : data = 13'b0000001101001;
			8'b01101010 : data = 13'b0000001101010;
			8'b01101011 : data = 13'b0000001101011;
			8'b01101100 : data = 13'b0000001101100;
			8'b01101101 : data = 13'b0000001101101;
			8'b01101110 : data = 13'b0000001101110;
			8'b01101111 : data = 13'b0000001101111;
			8'b01110000 : data = 13'b0000001110000;
			8'b01110001 : data = 13'b0000001110001;
			8'b01110010 : data = 13'b0000001110010;
			8'b01110011 : data = 13'b0000001110011;
			8'b01110100 : data = 13'b0000001110100;
			8'b01110101 : data = 13'b0000001110101;
			8'b01110110 : data = 13'b0000001110110;
			8'b01110111 : data = 13'b0000001110111;
			8'b01111000 : data = 13'b0000001111000;
			8'b01111001 : data = 13'b0000001111001;
			8'b01111010 : data = 13'b0000001111010;
			8'b01111011 : data = 13'b0000001111011;
			8'b01111100 : data = 13'b0000001111100;
			8'b01111101 : data = 13'b0000001111101;
			8'b01111110 : data = 13'b0000001111110;
			8'b01111111 : data = 13'b0000001111111;
			8'b10000000 : data = 13'b0000010000000;
			8'b10000001 : data = 13'b0000010000001;
			8'b10000010 : data = 13'b0000010000010;
			8'b10000011 : data = 13'b0000010000011;
			8'b10000100 : data = 13'b0000010000100;
			8'b10000101 : data = 13'b0000010000101;
			8'b10000110 : data = 13'b0000010000110;
			8'b10000111 : data = 13'b0000010000111;
			8'b10001000 : data = 13'b0000010001000;
			8'b10001001 : data = 13'b0000010001001;
			8'b10001010 : data = 13'b0000010001010;
			8'b10001011 : data = 13'b0000010001011;
			8'b10001100 : data = 13'b0000010001100;
			8'b10001101 : data = 13'b0000010001101;
			8'b10001110 : data = 13'b0000010001110;
			8'b10001111 : data = 13'b0000010001111;
			8'b10010000 : data = 13'b0000010010000;
			8'b10010001 : data = 13'b0000010010001;
			8'b10010010 : data = 13'b0000010010010;
			8'b10010011 : data = 13'b0000010010011;
			8'b10010100 : data = 13'b0000010010100;
			8'b10010101 : data = 13'b0000010010101;
			8'b10010110 : data = 13'b0000010010110;
			8'b10010111 : data = 13'b0000010010111;
			8'b10011000 : data = 13'b0000010011000;
			8'b10011001 : data = 13'b0000010011001;
			8'b10011010 : data = 13'b0000010011010;
			8'b10011011 : data = 13'b0000010011011;
			8'b10011100 : data = 13'b0000010011100;
			8'b10011101 : data = 13'b0000010011101;
			8'b10011110 : data = 13'b0000010011110;
			8'b10011111 : data = 13'b0000010011111;
			8'b10100000 : data = 13'b0000010100000;
			8'b10100001 : data = 13'b0000010100001;
			8'b10100010 : data = 13'b0000010100010;
			8'b10100011 : data = 13'b0000010100011;
			8'b10100100 : data = 13'b0000010100100;
			8'b10100101 : data = 13'b0000010100101;
			8'b10100110 : data = 13'b0000010100110;
			8'b10100111 : data = 13'b0000010100111;
			8'b10101000 : data = 13'b0000010101000;
			8'b10101001 : data = 13'b0000010101001;
			8'b10101010 : data = 13'b0000010101010;
			8'b10101011 : data = 13'b0000010101011;
			8'b10101100 : data = 13'b0000010101100;
			8'b10101101 : data = 13'b0000010101101;
			8'b10101110 : data = 13'b0000010101110;
			8'b10101111 : data = 13'b0000010101111;
			8'b10110000 : data = 13'b0000010110000;
			8'b10110001 : data = 13'b0000010110001;
			8'b10110010 : data = 13'b0000010110010;
			8'b10110011 : data = 13'b0000010110011;
			8'b10110100 : data = 13'b0000010110100;
			8'b10110101 : data = 13'b0000010110101;
			8'b10110110 : data = 13'b0000010110110;
			8'b10110111 : data = 13'b0000010110111;
			8'b10111000 : data = 13'b0000010111000;
			8'b10111001 : data = 13'b0000010111001;
			8'b10111010 : data = 13'b0000010111010;
			8'b10111011 : data = 13'b0000010111011;
			8'b10111100 : data = 13'b0000010111100;
			8'b10111101 : data = 13'b0000010111101;
			8'b10111110 : data = 13'b0000010111110;
			8'b10111111 : data = 13'b0000010111111;
			8'b11000000 : data = 13'b0000011000000;
			8'b11000001 : data = 13'b0000011000001;
			8'b11000010 : data = 13'b0000011000010;
			8'b11000011 : data = 13'b0000011000011;
			8'b11000100 : data = 13'b0000011000100;
			8'b11000101 : data = 13'b0000011000101;
			8'b11000110 : data = 13'b0000011000110;
			8'b11000111 : data = 13'b0000011000111;
			8'b11001000 : data = 13'b0000011001000;
			8'b11001001 : data = 13'b0000011001001;
			8'b11001010 : data = 13'b0000011001010;
			8'b11001011 : data = 13'b0000011001011;
			8'b11001100 : data = 13'b0000011001100;
			8'b11001101 : data = 13'b0000011001101;
			8'b11001110 : data = 13'b0000011001110;
			8'b11001111 : data = 13'b0000011001111;
			8'b11010000 : data = 13'b0000011010000;
			8'b11010001 : data = 13'b0000011010001;
			8'b11010010 : data = 13'b0000011010010;
			8'b11010011 : data = 13'b0000011010011;
			8'b11010100 : data = 13'b0000011010100;
			8'b11010101 : data = 13'b0000011010101;
			8'b11010110 : data = 13'b0000011010110;
			8'b11010111 : data = 13'b0000011010111;
			8'b11011000 : data = 13'b0000011011000;
			8'b11011001 : data = 13'b0000011011001;
			8'b11011010 : data = 13'b0000011011010;
			8'b11011011 : data = 13'b0000011011011;
			8'b11011100 : data = 13'b0000011011100;
			8'b11011101 : data = 13'b0000011011101;
			8'b11011110 : data = 13'b0000011011110;
			8'b11011111 : data = 13'b0000011011111;
			8'b11100000 : data = 13'b0000011100000;
			8'b11100001 : data = 13'b0000011100001;
			8'b11100010 : data = 13'b0000011100010;
			8'b11100011 : data = 13'b0000011100011;
			8'b11100100 : data = 13'b0000011100100;
			8'b11100101 : data = 13'b0000011100101;
			8'b11100110 : data = 13'b0000011100110;
			8'b11100111 : data = 13'b0000011100111;
			8'b11101000 : data = 13'b0000011101000;
			8'b11101001 : data = 13'b0000011101001;
			8'b11101010 : data = 13'b0000011101010;
			8'b11101011 : data = 13'b0000011101011;
			8'b11101100 : data = 13'b0000011101100;
			8'b11101101 : data = 13'b0000011101101;
			8'b11101110 : data = 13'b0000011101110;
			8'b11101111 : data = 13'b0000011101111;
			8'b11110000 : data = 13'b0000011110000;
			8'b11110001 : data = 13'b0000011110001;
			8'b11110010 : data = 13'b0000011110010;
			8'b11110011 : data = 13'b0000011110011;
			8'b11110100 : data = 13'b0000011110100;
			8'b11110101 : data = 13'b0000011110101;
			8'b11110110 : data = 13'b0000011110110;
			8'b11110111 : data = 13'b0000011110111;
			8'b11111000 : data = 13'b0000011111000;
			8'b11111001 : data = 13'b0000011111001;
			8'b11111010 : data = 13'b0000011111010;
			8'b11111011 : data = 13'b0000011111011;
			8'b11111100 : data = 13'b0000011111100;
			8'b11111101 : data = 13'b0000011111101;
			8'b11111110 : data = 13'b0000011111110;
			8'b11111111 : data = 13'b0000011111111;


         default : data = 8'b0000000000000; 
	 endcase
	 end
	
end    

endmodule 